`timescale 1ns/1ps

module alu_test;
reg [31:0] instruction, regA, regB;
wire [31:0] result;
wire [2:0] flags;
reg [31:0] correct_result;
ALU testalu(instruction, regA, regB, result, flags);
initial 
begin
$display("instruction:op:func:  regA  :  regB  :flags: result :correct_result");
$monitor("   %h:%h: %h :%h:%h: %b :%h:%h",
instruction, testalu.opcode, testalu.funct, regA, regB, flags, result, correct_result);
// add: 1 + 2
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_0000;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;

// add: overflow
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_0000;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1110;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_0001;
correct_result <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;

// addi: 1 + 2(imm)
#10 instruction <= 32'b0010_0000_0010_0010_0000_0000_0000_0010;
regA <= 32'b1;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;

// addi: 3 + -1(imm)
#10 instruction <= 32'b0010_0000_0010_0010_1111_1111_1111_1111;
regA <= 32'b0;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;

// addi: overflow
#10 instruction <= 32'b0010_0000_0010_0010_1111_1111_1111_1111;
regA <= 32'b0;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
correct_result <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;

// addu
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_0001;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

// addiu:
#10 instruction <= 32'b0010_0100_0000_0010_0000_0000_0000_0001;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b0;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

// sub:
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_0010;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;

// sub: overflow
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_0010;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
correct_result <= 32'b1000_0000_0000_0000_0000_0000_0000_0011;

// subu:
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_0011;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
correct_result <= 32'b0000_0000_0000_0000_0000_0000;

// and:
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_0100;
regA <= 32'b0000_0110_0000_0000_0000_1100_0000_1111;
regB <= 32'b0000_0110_0000_0000_0000_0110_0000_1110;
correct_result <= 32'b0000_0110_0000_1000_0000_0100_0000_1110;

// andi:
#10 instruction <= 32'b0011_0000_0010_0010_1111_1111_1111_1110;
regA <= 32'b0;
regB <= 32'b0000_0000_0000_0000_0000_1100_0000_0011;
correct_result <= 32'b0000_0000_0000_0000_0000_1100_0000_0010;

//nor:
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_0111;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b0000_0110_0000_1100_0000_0110_0000_0011;
correct_result <= 32'b0000_0000_0000_0000_0000_0000;

//or:
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_0101;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b0000_0110_0000_1100_0000_0110_0000_0011;
correct_result <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;

//ori:
#10 instruction <= 32'b0011_0100_0010_0010_1111_1111_1111_1110;
regA <= 32'b0;
regB <= 32'b0000_0000_0000_0000_0000_1100_0000_0010;
correct_result <= 32'b0000_0000_0000_0000_1111_1111_1111_1110;

//xor:
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_0110;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b0000_0110_0000_1100_0000_0110_0000_0011;
correct_result <= 32'b1111_1001_1111_0011_1111_1001_1111_1100;

//xori
#10 instruction <= 32'b0011_1000_0010_0010_1111_1111_1111_1111;
regA <= 32'b0;
regB <= 32'b0000_0000_0000_0000_0000_1100_0000_0011;
correct_result <= 32'b0000_0000_0000_0000_1111_0011_1111_1100;

//beq:
#10 instruction <= 32'b0001_0000_0000_0001_0000_0000_0000_0000;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

//beq:
#10 instruction <= 32'b0001_0000_0000_0001_0000_0000_0000_0000;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//bne equal
#10 instruction <= 32'b0001_0100_0000_0001_0000_0000_0000_0000;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//bne not equal
#10 instruction <= 32'b0001_0100_0000_0001_0000_0000_0000_0000;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
regB <= 32'b0000_0100_0110_1000_0000_1100_0000_0011;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

//slt bigger
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_1010;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
correct_result <= 32'b0;

//slt smaller
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_1010;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
regB <= 32'b0000_1100_0110_1000_0000_1100_0000_0011;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

//slti bigger
#10 instruction <= 32'b0010_1000_0000_0001_0000_0000_0000_0000;
regA <= 32'b0000_0100_0110_1000_0000_1100_0000_0011;
regB <= 32'b0;
correct_result <= 32'b0;

//slti smaller
#10 instruction <= 32'b0010_1000_0000_0001_0111_1111_1111_1111;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
regB <= 32'b0;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

//sltiu: bigger
#10 instruction <= 32'b0010_1100_0000_0001_0010_0000_1100_0011;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b0;
correct_result <= 32'b0;

//sltiu: smaller
#10 instruction <= 32'b0010_1100_0000_0001_1111_1111_1111_1111;
regA <= 32'b0000_0000_0000_0000_0000_1100_0000_0011;
regB <= 32'b0;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

//sltu: bigger
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_1011;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b0000_0000_0000_0000_0000_1100_0000_0011;
correct_result <= 32'b0;

//sltu: smaller
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0010_1011;
regA <= 32'b0000_0000_0000_0000_0000_1100_0000_0011;
regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
correct_result <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

//lw
#10 instruction <= 32'b1000_1100_0000_0001_0000_0000_0000_0001;
regA <= 32'b0000_0000_0000_0000_0000_1100_0000_0011;
regB <= 32'b0;
correct_result <= 32'b0000_0000_0000_0000_0000_1100_0000_0100;

//sw
#10 instruction <= 32'b1000_1100_0000_0001_0000_0000_0000_0001;
regA <= 32'b0000_0000_0000_0000_0000_1100_0000_0011;
regB <= 32'b0;
correct_result <= 32'b0000_0000_0000_0000_0000_1100_0000_0100;

//sll 
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0100_0000;
regA <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;
regB <= 32'b1101_1101_1101_1101_1101_1101_1101_1101;
correct_result <= 32'b1011_1011_1011_1011_1011_1011_1011_1010;

//sllv:
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0000_0100;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
correct_result <= 32'b1111_1111_1111_1111_1111_1111_1111_1110;

//srl
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_1000_0010;
regA <= 32'b0;
regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
correct_result <= 32'b0011_1111_1111_1111_1111_1111_1111_1111;

//srlv:
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0000_0110;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
correct_result <= 32'b0011_1111_1111_1111_1111_1111_1111_1111;

//sra: negative
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0100_0011;
regA <= 32'b0;
regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
correct_result <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;

//sra: positive
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0100_0011;
regA <= 32'b0;
regB <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;
correct_result <= 32'b0011_1111_1111_1111_1111_1111_1111_1111;

//srav: negtive
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0000_0111;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
correct_result <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;

// test srav (positive regB >>> regA[4:0])
#10 instruction <= 32'b0000_0000_0000_0001_0001_0000_0000_0111;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;
correct_result <= 32'b0011_1111_1111_1111_1111_1111_1111_1111;

#10 $finish;
end
endmodule